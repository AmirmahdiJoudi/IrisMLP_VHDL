LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE layer_pkg IS
        TYPE BUS_ARRAY IS ARRAY(NATURAL RANGE <>) OF STD_LOGIC_VECTOR;
END PACKAGE;