LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE ARR_TYPE IS
    TYPE ARR IS ARRAY (NATURAL RANGE <>) OF INTEGER;
    TYPE ARR_STD IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR (200-1 DOWNTO 0);
END PACKAGE ARR_TYPE;